`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/07/2024 03:00:35 PM
// Design Name: 
// Module Name: regfile
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module regfile(
    input [63:0] WriteData,
    input [4:0] rs1,
    input [4:0] rs2,
    input [4:0] rd,
    input RegWrite,
    input clk,
    input reset,
    output reg [63:0]ReadData1,
    output reg [63:0]ReadData2
    );
    
    reg [63:0]registers[31:0];
    
    integer i;
    initial
    begin
    
    for (i=0; i<64 ;i = i+1)
    begin
    registers[i] = 0;
    end
    
    end
    
    always @(posedge clk)
    begin
    if (RegWrite)
        begin registers[rd] <= WriteData; end
    end
    
    always @(*)
    begin
    if (reset)
    begin
    ReadData1 = 64'b0;
    ReadData2 = 64'b0;
    end
    
    else
    begin
    ReadData1 = registers[rs1];
    ReadData2 = registers[rs2];
    end
    end

//    always @(rs1 or rs2 or reset or registers)
//    begin
//    ReadData1 = registers[rs1];
//    ReadData2 = registers[rs2];
    
//    if (reset)
//    begin
//    ReadData1 = 0;
//    ReadData2 = 0;
//    end
//    end
    
//    always @(RegWrite&&clk)
//    begin
//    registers[rd] = WriteData;
//    end
    
endmodule


//    registers[0] = 64'b0000000000000000000000000000000000000000000000000000000000000000;
//    registers[1] = 64'b0000000000000000000000000000000000000000000000000000000000000001;
//    registers[2] = 64'b0000000000000000000000000000000000000000000000000000000000000010;
//    registers[3] = 64'b0000000000000000000000000000000000000000000000000000000000000011;
//    registers[4] = 64'b0000000000000000000000000000000000000000000000000000000000000100;
//    registers[5] = 64'b0000000000000000000000000000000000000000000000000000000000000101;
//    registers[6] = 64'b0000000000000000000000000000000000000000000000000000000000000110;
//    registers[7] = 64'b0000000000000000000000000000000000000000000000000000000000000111;
//    registers[8] = 64'b0000000000000000000000000000000000000000000000000000000000001000;
//    registers[9] = 64'b0000000000000000000000000000000000000000000000000000000000001001;
//    registers[10] = 64'b0000000000000000000000000000000000000000000000000000000000001010;
//    registers[11] = 64'b0000000000000000000000000000000000000000000000000000000000001011;
//    registers[12] = 64'b0000000000000000000000000000000000000000000000000000000000001100;
//    registers[13] = 64'b0000000000000000000000000000000000000000000000000000000000001101;
//    registers[14] = 64'b0000000000000000000000000000000000000000000000000000000000001100;
//    registers[15] = 64'b0000000000000000000000000000000000000000000000000000000000001101;
//    registers[16] = 64'b0000000000000000000000000000000000000000000000000000000000010000;
//    registers[17] = 64'b0000000000000000000000000000000000000000000000000000000000010001;
//    registers[18] = 64'b0000000000000000000000000000000000000000000000000000000000010000;
//    registers[19] = 64'b0000000000000000000000000000000000000000000000000000000000010001;
//    registers[20] = 64'b0000000000000000000000000000000000000000000000000000000000010100;
//    registers[21] = 64'b0000000000000000000000000000000000000000000000000000000000010101;
//    registers[22] = 64'b0000000000000000000000000000000000000000000000000000000000010100;
//    registers[23] = 64'b0000000000000000000000000000000000000000000000000000000000010101;
//    registers[24] = 64'b0000000000000000000000000000000000000000000000000000000000011000;
//    registers[25] = 64'b0000000000000000000000000000000000000000000000000000000000011001;
//    registers[26] = 64'b0000000000000000000000000000000000000000000000000000000000011000;
//    registers[27] = 64'b0000000000000000000000000000000000000000000000000000000000011001;
//    registers[28] = 64'b0000000000000000000000000000000000000000000000000000000000011100;
//    registers[29] = 64'b0000000000000000000000000000000000000000000000000000000000011101;
//    registers[30] = 64'b0000000000000000000000000000000000000000000000000000000000011100;
//    registers[31] = 64'b0000000000000000000000000000000000000000000000000000000000011101;
